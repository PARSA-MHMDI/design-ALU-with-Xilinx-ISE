library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity decoder_3to8 is
	Port( a 	: in std_logic_vector(2 downto 0);
			q : out std_logic_vector(7 downto 0)
		  );
end decoder_3to8;

architecture Behavioral of decoder_3to8 is

begin

	with a select 
			q  <= "00000001" after 1 ns when "000" ,
					"00000010" after 1 ns when "001",
					"00000100" after 1 ns when "010",
					"00001000" after 1 ns when "011",
					"00010000" after 1 ns when "100",
					"00100000" after 1 ns when "101",
					"01000000" after 1 ns when "110",
					"10000000" after 1 ns when "111",

					"00000000" when others;
end Behavioral;

